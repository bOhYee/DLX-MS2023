LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE WORK.Globals.ALL;

ENTITY ND_GENERIC IS
	GENERIC(NBIT: integer := NumBit);

	PORT(A, B: IN std_logic_vector(NBIT-1 DOWNTO 0);
		 Y: OUT std_logic_vector(NBIT-1 DOWNTO 0));
END ND_GENERIC;


ARCHITECTURE BEHAVIOURAL OF ND_GENERIC IS
BEGIN

	AndProc: PROCESS(A,B)
	BEGIN
		Y <= NOT(A AND B);
	END PROCESS AndProc;

END BEHAVIOURAL;