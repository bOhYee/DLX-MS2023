LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE WORK.Globals.ALL;

ENTITY AND2_GENERIC IS
	GENERIC(NBIT: integer := NumBit);

	PORT(A, B:	IN std_logic_vector(NBIT-1 DOWNTO 0);
		 Y:	OUT	std_logic_vector(NBIT-1 DOWNTO 0));
END AND2_GENERIC;


ARCHITECTURE BEHAVIORAL of AND2_GENERIC IS
BEGIN

	AndProc: PROCESS(A, B)
	BEGIN
		Y <= A AND B;
	END PROCESS AndProc;

END BEHAVIORAL;