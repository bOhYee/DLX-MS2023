LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE WORK.Globals.ALL;

ENTITY PG_NETWORK is 
	PORT(A, B : IN std_logic;
		 P, G : OUT std_logic);	
END PG_NETWORK;

ARCHITECTURE BEHAVIORAL OF PG_NETWORK IS
BEGIN

	P <= A XOR B;
	G <= A AND B;

END BEHAVIORAL;