LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY GENERATE_BLOCK is 
	PORT(Ph, Gh, Gl: IN std_logic;
	     Ghl : OUT std_logic);	
END GENERATE_BLOCK;

ARCHITECTURE BEHAVIORAL OF GENERATE_BLOCK IS
BEGIN

	Ghl <= Gh OR (Ph AND Gl);
	
END BEHAVIORAL;
