LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE WORK.Globals.ALL;

ENTITY XOR2_GENERIC IS
	GENERIC(NBIT: integer := NumBit);

	PORT(A, B:	IN std_logic_vector(NBIT-1 DOWNTO 0);
		 Y:	OUT	std_logic_vector(NBIT-1 DOWNTO 0));
END XOR2_GENERIC;

ARCHITECTURE BEHAVIORAL of XOR2_GENERIC IS
BEGIN

	Xor2Proc: PROCESS(A, B)
	BEGIN
		Y <= A XOR B;
	END PROCESS Xor2Proc;

END BEHAVIORAL;