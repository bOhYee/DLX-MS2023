LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE WORK.Globals.ALL;

ENTITY IV_GENERIC IS
	GENERIC(NBIT: integer := NumBit);

	PORT(A:	IN std_logic_vector(NBIT-1 DOWNTO 0);
		 Y:	OUT	std_logic_vector(NBIT-1 DOWNTO 0));
END IV_GENERIC;


ARCHITECTURE BEHAVIORAL of IV_GENERIC IS
BEGIN

	InvProc: PROCESS(A)
	BEGIN
		Y <= NOT(A);
	END PROCESS InvProc;

END BEHAVIORAL;
