LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE WORK.Globals.ALL;

ENTITY OR2_GENERIC IS
	GENERIC(NBIT: integer := NumBit);

	PORT(A, B:	IN std_logic_vector(NBIT-1 DOWNTO 0);
		 Y:	OUT	std_logic_vector(NBIT-1 DOWNTO 0));
END OR2_GENERIC;

ARCHITECTURE BEHAVIORAL of OR2_GENERIC IS
BEGIN

	OrProc: PROCESS(A, B)
	BEGIN
		Y <= A OR B;
	END PROCESS OrProc;

END BEHAVIORAL;
